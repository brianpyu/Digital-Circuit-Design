// processor.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module processor (
		output wire [10:0] address_external_connection_export,           //           address_external_connection.export
		input  wire        characterreceived_external_connection_export, // characterreceived_external_connection.export
		input  wire        charactersent_external_connection_export,     //     charactersent_external_connection.export
		input  wire        clk_clk,                                      //                                   clk.clk
		inout  wire [7:0]  data_external_connection_export,              //              data_external_connection.export
		output wire        load_external_connection_export,              //              load_external_connection.export
		output wire        outputenable_external_connection_export,      //      outputenable_external_connection.export
		input  wire [7:0]  parallelinput_external_connection_export,     //     parallelinput_external_connection.export
		output wire [7:0]  paralleloutput_external_connection_export,    //    paralleloutput_external_connection.export
		input  wire        reset_reset_n,                                //                                 reset.reset_n
		output wire        transmitenable_external_connection_export,    //    transmitenable_external_connection.export
		output wire        writeenable_external_connection_export        //       writeenable_external_connection.export
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [18:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [18:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_mem_s1_chipselect;                // mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	wire  [31:0] mm_interconnect_0_onchip_mem_s1_readdata;                  // onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_mem_s1_address;                   // mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	wire   [3:0] mm_interconnect_0_onchip_mem_s1_byteenable;                // mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	wire         mm_interconnect_0_onchip_mem_s1_write;                     // mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	wire  [31:0] mm_interconnect_0_onchip_mem_s1_writedata;                 // mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	wire         mm_interconnect_0_onchip_mem_s1_clken;                     // mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;             // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;               // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                  // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;              // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_paralleloutput_s1_chipselect;            // mm_interconnect_0:parallelOutput_s1_chipselect -> parallelOutput:chipselect
	wire  [31:0] mm_interconnect_0_paralleloutput_s1_readdata;              // parallelOutput:readdata -> mm_interconnect_0:parallelOutput_s1_readdata
	wire   [1:0] mm_interconnect_0_paralleloutput_s1_address;               // mm_interconnect_0:parallelOutput_s1_address -> parallelOutput:address
	wire         mm_interconnect_0_paralleloutput_s1_write;                 // mm_interconnect_0:parallelOutput_s1_write -> parallelOutput:write_n
	wire  [31:0] mm_interconnect_0_paralleloutput_s1_writedata;             // mm_interconnect_0:parallelOutput_s1_writedata -> parallelOutput:writedata
	wire  [31:0] mm_interconnect_0_parallelinput_s1_readdata;               // parallelInput:readdata -> mm_interconnect_0:parallelInput_s1_readdata
	wire   [1:0] mm_interconnect_0_parallelinput_s1_address;                // mm_interconnect_0:parallelInput_s1_address -> parallelInput:address
	wire         mm_interconnect_0_transmitenable_s1_chipselect;            // mm_interconnect_0:transmitEnable_s1_chipselect -> transmitEnable:chipselect
	wire  [31:0] mm_interconnect_0_transmitenable_s1_readdata;              // transmitEnable:readdata -> mm_interconnect_0:transmitEnable_s1_readdata
	wire   [1:0] mm_interconnect_0_transmitenable_s1_address;               // mm_interconnect_0:transmitEnable_s1_address -> transmitEnable:address
	wire         mm_interconnect_0_transmitenable_s1_write;                 // mm_interconnect_0:transmitEnable_s1_write -> transmitEnable:write_n
	wire  [31:0] mm_interconnect_0_transmitenable_s1_writedata;             // mm_interconnect_0:transmitEnable_s1_writedata -> transmitEnable:writedata
	wire         mm_interconnect_0_load_s1_chipselect;                      // mm_interconnect_0:load_s1_chipselect -> load:chipselect
	wire  [31:0] mm_interconnect_0_load_s1_readdata;                        // load:readdata -> mm_interconnect_0:load_s1_readdata
	wire   [1:0] mm_interconnect_0_load_s1_address;                         // mm_interconnect_0:load_s1_address -> load:address
	wire         mm_interconnect_0_load_s1_write;                           // mm_interconnect_0:load_s1_write -> load:write_n
	wire  [31:0] mm_interconnect_0_load_s1_writedata;                       // mm_interconnect_0:load_s1_writedata -> load:writedata
	wire  [31:0] mm_interconnect_0_characterreceived_s1_readdata;           // characterReceived:readdata -> mm_interconnect_0:characterReceived_s1_readdata
	wire   [1:0] mm_interconnect_0_characterreceived_s1_address;            // mm_interconnect_0:characterReceived_s1_address -> characterReceived:address
	wire  [31:0] mm_interconnect_0_charactersent_s1_readdata;               // characterSent:readdata -> mm_interconnect_0:characterSent_s1_readdata
	wire   [1:0] mm_interconnect_0_charactersent_s1_address;                // mm_interconnect_0:characterSent_s1_address -> characterSent:address
	wire         mm_interconnect_0_address_s1_chipselect;                   // mm_interconnect_0:address_s1_chipselect -> address:chipselect
	wire  [31:0] mm_interconnect_0_address_s1_readdata;                     // address:readdata -> mm_interconnect_0:address_s1_readdata
	wire   [1:0] mm_interconnect_0_address_s1_address;                      // mm_interconnect_0:address_s1_address -> address:address
	wire         mm_interconnect_0_address_s1_write;                        // mm_interconnect_0:address_s1_write -> address:write_n
	wire  [31:0] mm_interconnect_0_address_s1_writedata;                    // mm_interconnect_0:address_s1_writedata -> address:writedata
	wire         mm_interconnect_0_data_s1_chipselect;                      // mm_interconnect_0:data_s1_chipselect -> data:chipselect
	wire  [31:0] mm_interconnect_0_data_s1_readdata;                        // data:readdata -> mm_interconnect_0:data_s1_readdata
	wire   [1:0] mm_interconnect_0_data_s1_address;                         // mm_interconnect_0:data_s1_address -> data:address
	wire         mm_interconnect_0_data_s1_write;                           // mm_interconnect_0:data_s1_write -> data:write_n
	wire  [31:0] mm_interconnect_0_data_s1_writedata;                       // mm_interconnect_0:data_s1_writedata -> data:writedata
	wire         mm_interconnect_0_outputenable_s1_chipselect;              // mm_interconnect_0:outputEnable_s1_chipselect -> outputEnable:chipselect
	wire  [31:0] mm_interconnect_0_outputenable_s1_readdata;                // outputEnable:readdata -> mm_interconnect_0:outputEnable_s1_readdata
	wire   [1:0] mm_interconnect_0_outputenable_s1_address;                 // mm_interconnect_0:outputEnable_s1_address -> outputEnable:address
	wire         mm_interconnect_0_outputenable_s1_write;                   // mm_interconnect_0:outputEnable_s1_write -> outputEnable:write_n
	wire  [31:0] mm_interconnect_0_outputenable_s1_writedata;               // mm_interconnect_0:outputEnable_s1_writedata -> outputEnable:writedata
	wire         mm_interconnect_0_writeenable_s1_chipselect;               // mm_interconnect_0:writeEnable_s1_chipselect -> writeEnable:chipselect
	wire  [31:0] mm_interconnect_0_writeenable_s1_readdata;                 // writeEnable:readdata -> mm_interconnect_0:writeEnable_s1_readdata
	wire   [1:0] mm_interconnect_0_writeenable_s1_address;                  // mm_interconnect_0:writeEnable_s1_address -> writeEnable:address
	wire         mm_interconnect_0_writeenable_s1_write;                    // mm_interconnect_0:writeEnable_s1_write -> writeEnable:write_n
	wire  [31:0] mm_interconnect_0_writeenable_s1_writedata;                // mm_interconnect_0:writeEnable_s1_writedata -> writeEnable:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // sys_clk_timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [address:reset_n, characterReceived:reset_n, characterSent:reset_n, cpu:reset_n, data:reset_n, irq_mapper:reset, jtag_uart:rst_n, load:reset_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_mem:reset, outputEnable:reset_n, parallelInput:reset_n, parallelOutput:reset_n, rst_translator:in_reset, sys_clk_timer:reset_n, sysid:reset_n, transmitEnable:reset_n, writeEnable:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]

	processor_address address (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_address_s1_readdata),   //                    .readdata
		.out_port   (address_external_connection_export)       // external_connection.export
	);

	processor_characterReceived characterreceived (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_characterreceived_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_characterreceived_s1_readdata), //                    .readdata
		.in_port  (characterreceived_external_connection_export)     // external_connection.export
	);

	processor_characterReceived charactersent (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_charactersent_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_charactersent_s1_readdata), //                    .readdata
		.in_port  (charactersent_external_connection_export)     // external_connection.export
	);

	processor_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                    //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	processor_data data (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_s1_readdata),   //                    .readdata
		.bidir_port (data_external_connection_export)       // external_connection.export
	);

	processor_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	processor_load load (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_load_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_load_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_load_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_load_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_load_s1_readdata),   //                    .readdata
		.out_port   (load_external_connection_export)       // external_connection.export
	);

	processor_onchip_mem onchip_mem (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	processor_load outputenable (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_outputenable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_outputenable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_outputenable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_outputenable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_outputenable_s1_readdata),   //                    .readdata
		.out_port   (outputenable_external_connection_export)       // external_connection.export
	);

	processor_parallelInput parallelinput (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_parallelinput_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_parallelinput_s1_readdata), //                    .readdata
		.in_port  (parallelinput_external_connection_export)     // external_connection.export
	);

	processor_parallelOutput paralleloutput (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_paralleloutput_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_paralleloutput_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_paralleloutput_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_paralleloutput_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_paralleloutput_s1_readdata),   //                    .readdata
		.out_port   (paralleloutput_external_connection_export)       // external_connection.export
	);

	processor_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                       //   irq.irq
	);

	processor_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	processor_load transmitenable (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_transmitenable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmitenable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmitenable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmitenable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmitenable_s1_readdata),   //                    .readdata
		.out_port   (transmitenable_external_connection_export)       // external_connection.export
	);

	processor_load writeenable (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_writeenable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_writeenable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_writeenable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_writeenable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_writeenable_s1_readdata),   //                    .readdata
		.out_port   (writeenable_external_connection_export)       // external_connection.export
	);

	processor_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                                   //                         clk_0_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                   cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                  .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                  .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                  .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                  .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                  .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                  .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                  .readdata
		.cpu_instruction_master_readdatavalid    (cpu_instruction_master_readdatavalid),                      //                                  .readdatavalid
		.address_s1_address                      (mm_interconnect_0_address_s1_address),                      //                        address_s1.address
		.address_s1_write                        (mm_interconnect_0_address_s1_write),                        //                                  .write
		.address_s1_readdata                     (mm_interconnect_0_address_s1_readdata),                     //                                  .readdata
		.address_s1_writedata                    (mm_interconnect_0_address_s1_writedata),                    //                                  .writedata
		.address_s1_chipselect                   (mm_interconnect_0_address_s1_chipselect),                   //                                  .chipselect
		.characterReceived_s1_address            (mm_interconnect_0_characterreceived_s1_address),            //              characterReceived_s1.address
		.characterReceived_s1_readdata           (mm_interconnect_0_characterreceived_s1_readdata),           //                                  .readdata
		.characterSent_s1_address                (mm_interconnect_0_charactersent_s1_address),                //                  characterSent_s1.address
		.characterSent_s1_readdata               (mm_interconnect_0_charactersent_s1_readdata),               //                                  .readdata
		.cpu_jtag_debug_module_address           (mm_interconnect_0_cpu_jtag_debug_module_address),           //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write             (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                  .write
		.cpu_jtag_debug_module_read              (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                  .read
		.cpu_jtag_debug_module_readdata          (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                  .readdata
		.cpu_jtag_debug_module_writedata         (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                  .writedata
		.cpu_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                  .debugaccess
		.data_s1_address                         (mm_interconnect_0_data_s1_address),                         //                           data_s1.address
		.data_s1_write                           (mm_interconnect_0_data_s1_write),                           //                                  .write
		.data_s1_readdata                        (mm_interconnect_0_data_s1_readdata),                        //                                  .readdata
		.data_s1_writedata                       (mm_interconnect_0_data_s1_writedata),                       //                                  .writedata
		.data_s1_chipselect                      (mm_interconnect_0_data_s1_chipselect),                      //                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.load_s1_address                         (mm_interconnect_0_load_s1_address),                         //                           load_s1.address
		.load_s1_write                           (mm_interconnect_0_load_s1_write),                           //                                  .write
		.load_s1_readdata                        (mm_interconnect_0_load_s1_readdata),                        //                                  .readdata
		.load_s1_writedata                       (mm_interconnect_0_load_s1_writedata),                       //                                  .writedata
		.load_s1_chipselect                      (mm_interconnect_0_load_s1_chipselect),                      //                                  .chipselect
		.onchip_mem_s1_address                   (mm_interconnect_0_onchip_mem_s1_address),                   //                     onchip_mem_s1.address
		.onchip_mem_s1_write                     (mm_interconnect_0_onchip_mem_s1_write),                     //                                  .write
		.onchip_mem_s1_readdata                  (mm_interconnect_0_onchip_mem_s1_readdata),                  //                                  .readdata
		.onchip_mem_s1_writedata                 (mm_interconnect_0_onchip_mem_s1_writedata),                 //                                  .writedata
		.onchip_mem_s1_byteenable                (mm_interconnect_0_onchip_mem_s1_byteenable),                //                                  .byteenable
		.onchip_mem_s1_chipselect                (mm_interconnect_0_onchip_mem_s1_chipselect),                //                                  .chipselect
		.onchip_mem_s1_clken                     (mm_interconnect_0_onchip_mem_s1_clken),                     //                                  .clken
		.outputEnable_s1_address                 (mm_interconnect_0_outputenable_s1_address),                 //                   outputEnable_s1.address
		.outputEnable_s1_write                   (mm_interconnect_0_outputenable_s1_write),                   //                                  .write
		.outputEnable_s1_readdata                (mm_interconnect_0_outputenable_s1_readdata),                //                                  .readdata
		.outputEnable_s1_writedata               (mm_interconnect_0_outputenable_s1_writedata),               //                                  .writedata
		.outputEnable_s1_chipselect              (mm_interconnect_0_outputenable_s1_chipselect),              //                                  .chipselect
		.parallelInput_s1_address                (mm_interconnect_0_parallelinput_s1_address),                //                  parallelInput_s1.address
		.parallelInput_s1_readdata               (mm_interconnect_0_parallelinput_s1_readdata),               //                                  .readdata
		.parallelOutput_s1_address               (mm_interconnect_0_paralleloutput_s1_address),               //                 parallelOutput_s1.address
		.parallelOutput_s1_write                 (mm_interconnect_0_paralleloutput_s1_write),                 //                                  .write
		.parallelOutput_s1_readdata              (mm_interconnect_0_paralleloutput_s1_readdata),              //                                  .readdata
		.parallelOutput_s1_writedata             (mm_interconnect_0_paralleloutput_s1_writedata),             //                                  .writedata
		.parallelOutput_s1_chipselect            (mm_interconnect_0_paralleloutput_s1_chipselect),            //                                  .chipselect
		.sys_clk_timer_s1_address                (mm_interconnect_0_sys_clk_timer_s1_address),                //                  sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                  (mm_interconnect_0_sys_clk_timer_s1_write),                  //                                  .write
		.sys_clk_timer_s1_readdata               (mm_interconnect_0_sys_clk_timer_s1_readdata),               //                                  .readdata
		.sys_clk_timer_s1_writedata              (mm_interconnect_0_sys_clk_timer_s1_writedata),              //                                  .writedata
		.sys_clk_timer_s1_chipselect             (mm_interconnect_0_sys_clk_timer_s1_chipselect),             //                                  .chipselect
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //               sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),            //                                  .readdata
		.transmitEnable_s1_address               (mm_interconnect_0_transmitenable_s1_address),               //                 transmitEnable_s1.address
		.transmitEnable_s1_write                 (mm_interconnect_0_transmitenable_s1_write),                 //                                  .write
		.transmitEnable_s1_readdata              (mm_interconnect_0_transmitenable_s1_readdata),              //                                  .readdata
		.transmitEnable_s1_writedata             (mm_interconnect_0_transmitenable_s1_writedata),             //                                  .writedata
		.transmitEnable_s1_chipselect            (mm_interconnect_0_transmitenable_s1_chipselect),            //                                  .chipselect
		.writeEnable_s1_address                  (mm_interconnect_0_writeenable_s1_address),                  //                    writeEnable_s1.address
		.writeEnable_s1_write                    (mm_interconnect_0_writeenable_s1_write),                    //                                  .write
		.writeEnable_s1_readdata                 (mm_interconnect_0_writeenable_s1_readdata),                 //                                  .readdata
		.writeEnable_s1_writedata                (mm_interconnect_0_writeenable_s1_writedata),                //                                  .writedata
		.writeEnable_s1_chipselect               (mm_interconnect_0_writeenable_s1_chipselect)                //                                  .chipselect
	);

	processor_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
